`include "src/modules/serial_com.sv"